library verilog;
use verilog.vl_types.all;
entity GCD_vlg_vec_tst is
end GCD_vlg_vec_tst;
